// code to be simplified 

class 
